module rx (
    input clk,
    input rst,
    input rx,

    output reg rx_bit,
    output reg rx_bit_rdy
);
    
endmodule